module overflow(a, b, out);
	input[31:0] a,b;
	output out;
	
	

endmodule
